root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1142.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1143.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1144.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1145.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1146.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1147.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1148.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1149.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1150.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1151.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1152.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1153.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1154.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1155.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1156.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1157.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1158.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1159.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1160.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1161.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1162.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1163.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1164.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1165.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1166.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1167.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1168.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1169.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1170.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1171.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1172.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1173.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1174.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1175.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1176.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1177.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1178.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1179.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1180.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0001/stopFlatNtuples_1181.root
