root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3640.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3641.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3642.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3643.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3644.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3645.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3646.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3647.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3648.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3649.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3650.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3651.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3652.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3653.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3654.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3655.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3656.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3657.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3658.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3659.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3660.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3661.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3662.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3663.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3664.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3665.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3666.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3667.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3668.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3669.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3670.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3671.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3672.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3673.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3674.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3675.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3676.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3677.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3678.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0003/stopFlatNtuples_3679.root
