root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3702.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3703.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3704.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3705.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3706.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3707.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3708.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3709.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3710.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3711.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3712.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3713.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3714.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3715.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3716.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3717.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3718.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3719.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3720.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3721.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3722.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3723.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3724.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3725.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3726.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3727.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3728.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3729.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3730.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3731.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3732.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3733.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3734.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3735.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3736.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3737.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3738.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3739.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3740.root
root://cmseos.fnal.gov//store/user/lpcsusyhad/Stop_production/Spring16_80X_Nov_2016_Ntp_v11X_new_IDs/MET/Spring16_80X_Nov_2016_Ntp_v11p0_new_IDs_MET-Run2016H-PromptReco-v2/161111_231134/0003/stopFlatNtuples_3741.root
