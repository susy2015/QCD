root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1080.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1081.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1082.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1083.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1084.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1085.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1086.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1087.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1088.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1089.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1090.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1091.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1092.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1093.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1094.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1095.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1096.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1097.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1098.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1099.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1100.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1101.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1102.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1103.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1104.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1105.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1106.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1107.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1108.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1109.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1110.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1111.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1112.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1113.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1114.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1115.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1116.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1117.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1118.root
root://cmseos.fnal.gov//store/group/lpcsusyhad/Stop_production/Summer16_80X_Jan_2017_Ntp_v12X/MET/Summer16_80X_Jan_2017_Ntp_v12p0_MET-Run2016H-PromptReco-v2/170126_214332/0001/stopFlatNtuples_1119.root
